Library IEEE;
Use IEEE.Std_logic_1164.all;


Entity Coefficients_A is
	PORT(
	SEL : in Std_logic_vector(3 downto 0);
	QOUT: out Std_logic_vector(63 downto 0)
	
	);
End Entity Coefficients_A; 

Architecture DataFlow of Coefficients_A is
Begin	
	
OROM_A : process(SEL)    
begin  
    case SEL is
        when "0000" => QOUT <= "0000000000000001000000000000000000000000000000000000000000000000";
        when "0001" => QOUT <= "1111111111111110010100111001110010011001111100000100101010101100";
        when "0010" => QOUT <= "1111111111111101100010010010100010001100000111110010001001111010";
        when "0011" => QOUT <= "0000000000000011100101010110110100000000101111111011000011110000";
        when "0100" => QOUT <= "0000000000000101000010011101110100100010000101010001011111110011";
        when "0101" => QOUT <= "1111111111111011001111011011010001101000111101100101010111011111";
        when "0110" => QOUT <= "1111111111111010100111101010100001110011111111010010010001110111";
        when "0111" => QOUT <= "0000000000000010110000111011110000010101001010111010100010000000";
        when "1000" => QOUT <= "0000000000000100000010000001011011100000000010100110101111110100";
        when "1001" => QOUT <= "1111111111111111000001110011100000111000001101101111011001001011";
        when "1010" => QOUT <= "1111111111111110100011101000011110101100100111110100010100100000";
        when "1011" => QOUT <= "1111111111111111111011110101000001100100010010001001101110101100";
        when "1100" => QOUT <= "0000000000000000010101101011000010011100010101100101010101110011";
        when others => QOUT <= (others => '0');
    end case; 
end process OROM_A;

End Architecture DataFlow;


 
