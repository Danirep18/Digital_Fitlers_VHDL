Library IEEE;
Use IEEE.Std_logic_1164.all;


Entity Coefficients_B is
	PORT(
	SEL : in Std_logic_vector(3 downto 0);
	QOUT: out Std_logic_vector(63 downto 0)
	
	);
End Entity Coefficients_B; 

Architecture DataFlow of Coefficients_B is
Begin	
	
OROM_A : process(SEL)    
begin  
    case SEL is
        when "0000" => QOUT <= "0000000000000000011101101110000011010100000101101111001010111001";
        when "0001" => QOUT <= "1111111111111111110001010101001101011000001101111011010101100000";
        when "0010" => QOUT <= "1111111111111101101101010000011011011101111000011001000101111111";
        when "0011" => QOUT <= "0000000000000000100011100000100110101111100000001001001001111011";
        when "0100" => QOUT <= "0000000000000101010000110001100000111110000111110001110010110010";
        when "0101" => QOUT <= "1111111111111111101010000001100101010001011111110000100111101000";
        when "0110" => QOUT <= "1111111111111001001010110001001101101101011001100011111010101111";
        when "0111" => QOUT <= "1111111111111111101010000001100101010001011111110000100111101000";
        when "1000" => QOUT <= "0000000000000101010000110001100000111110000111110001110010110010";
        when "1001" => QOUT <= "0000000000000000100011100000100110101111100000001001001001111101";
        when "1010" => QOUT <= "1111111111111101101101010000011011011101111000011001000101111110";
        when "1011" => QOUT <= "1111111111111111110001010101001101011000001101111011010101100000";
        when "1100" => QOUT <= "0000000000000000011101101110000011010100000101101111001010111010";
        when others => QOUT <= (others => '0');
    end case; 
end process OROM_A;

End Architecture DataFlow;


 
